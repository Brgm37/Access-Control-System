library ieee;
use ieee.std_logic_1164.all;

	entity RingBuffer_tb is
	end RingBuffer_tb;
	
architecture RingBuffer_tb_arch of RingBuffer_tb is

	component RingBuffer is
		port(
			D: in std_logic_vector(3 downto 0);
			Q: out std_logic_vector(3 downto 0);
			CTS: in std_logic;
			clk: in std_logic;
			rst: in std_logic;
			DAV: in std_logic;
			Wreg: out std_logic;
			DAC: out std_logic
		); 
	end component;
	
	constant MCLK_PERIOD : time := 20 ns;
	constant MCLK_HALF_PERIOD : time := MCLK_PERIOD / 2;
	
	signal Dav_tb, CTS_tb, clk_tb, rst_tb, Wreg_tb, Dac_tb: std_logic;
	signal D_tb, Q_tb: std_logic_vector(3 downto 0);
	
	begin 
	
-- unit under Test 
	
	UUT: RingBuffer
		port map (
			D => D_tb,
			Q => Q_tb,
			CTS => CTS_tb,
			clk => clk_tb,
			rst => rst_tb,
			DAV => Dav_tb,
			Wreg => Wreg_tb,
			DAC => Dac_tb
		); 
	

	clk_gen : process
	begin
		clk_tb <= '0';
		wait for MCLK_HALF_PERIOD; 
		clk_tb <= '1';
		wait for MCLK_HALF_PERIOD;
	end process;
	
	
	-- 400 ns necessary to complete the test bench
	stimulus: process 
	begin
	
		-- reset
		rst_tb <= '1';
		dav_tb <= '0';
		cts_tb <= '0';
		wait for MCLK_PERIOD*2;
		
		rst_tb <= '0';
		
		wait for MCLK_PERIOD*2;
		
		cts_tb <= '1';
		
		wait for MCLK_PERIOD*2;
		
		dav_tb <= '1';
		D_tb <= "1111";
		
		wait for MCLK_PERIOD*2;
		
		
		wait for MCLK_PERIOD*2;
		
		
		wait for MCLK_PERIOD*2;
		
		
		dav_tb <= '0';
		
		wait for MCLK_PERIOD*2;
		
		cts_tb <= '1';
		
		wait for MCLK_PERIOD*6;
		
		--expecting Wreg == '1'
		-- expcting Q_tb == "1111"
		
		CTS_tb <= '0';
		
		wait for MCLK_PERIOD*2;
		
		
		D_tb <= "1010";
		dav_tb <= '1';
		
		wait for MCLK_PERIOD*2;
		
		
		wait for MCLK_PERIOD*2;
		
		
		wait for MCLK_PERIOD*2;
		
		
		dav_tb <= '0';
		
		wait for MCLK_PERIOD*2;
		
		D_tb <= "1011";
		dav_tb <= '1';
		
		wait for MCLK_PERIOD*2;
		
		
		wait for MCLK_PERIOD*2;
		
		
		wait for MCLK_PERIOD*2;
		
		
		dav_tb <= '0';
		
		wait for MCLK_PERIOD*2;
		
		cts_tb <= '1';
		
		wait for MCLK_PERIOD*6;
		
		--expecting Wreg == '1'
		-- expcting Q_tb == "1010"
		
		cts_tb <= '0';
		
		wait for MCLK_PERIOD*2;
		
		cts_tb <= '1';
		
		wait for MCLK_PERIOD*6;
		
		--expecting Wreg == '1'
		-- expcting Q_tb == "1011"
		
		CTS_tb <= '0';
		
		wait;
	end process;


end RingBuffer_tb_arch;